module head

pub fn head<T>(ls []T) T {
	return ls[0]
}