module vhs

