module vhs

fn main() {
	println('hi')
}
